--hello world file