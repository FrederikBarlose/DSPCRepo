-- CPU_System.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity CPU_System is
	port (
		clk_50                                    : in    std_logic                     := '0';             --                    clk_50_clk_in.clk
		dram_addr                                 : out   std_logic_vector(12 downto 0);                    --                             dram.addr
		dram_ba                                   : out   std_logic_vector(1 downto 0);                     --                                 .ba
		dram_cas_n                                : out   std_logic;                                        --                                 .cas_n
		dram_cke                                  : out   std_logic;                                        --                                 .cke
		dram_cs_n                                 : out   std_logic;                                        --                                 .cs_n
		dram_dq                                   : inout std_logic_vector(15 downto 0) := (others => '0'); --                                 .dq
		dram_dqm                                  : out   std_logic_vector(1 downto 0);                     --                                 .dqm
		dram_ras_n                                : out   std_logic;                                        --                                 .ras_n
		dram_we_n                                 : out   std_logic;                                        --                                 .we_n
		dram_clk_clk                              : out   std_logic;                                        --                         dram_clk.clk
		jtag_uart_0_avalon_jtag_slave_chipselect  : in    std_logic                     := '0';             --    jtag_uart_0_avalon_jtag_slave.chipselect
		jtag_uart_0_avalon_jtag_slave_address     : in    std_logic                     := '0';             --                                 .address
		jtag_uart_0_avalon_jtag_slave_read_n      : in    std_logic                     := '0';             --                                 .read_n
		jtag_uart_0_avalon_jtag_slave_readdata    : out   std_logic_vector(31 downto 0);                    --                                 .readdata
		jtag_uart_0_avalon_jtag_slave_write_n     : in    std_logic                     := '0';             --                                 .write_n
		jtag_uart_0_avalon_jtag_slave_writedata   : in    std_logic_vector(31 downto 0) := (others => '0'); --                                 .writedata
		jtag_uart_0_avalon_jtag_slave_waitrequest : out   std_logic;                                        --                                 .waitrequest
		in_port_to_the_pio_input_0                : in    std_logic_vector(7 downto 0)  := (others => '0'); --  pio_input_0_external_connection.export
		out_port_from_the_pio_output_0            : out   std_logic_vector(7 downto 0);                     -- pio_output_0_external_connection.export
		reset_reset_n                             : in    std_logic                     := '0'              --                            reset.reset_n
	);
end entity CPU_System;

architecture rtl of CPU_System is
	component mm_bus_counter is
		port (
			csi_clockreset_clk     : in  std_logic                     := 'X';             -- clk
			csi_clockreset_reset_n : in  std_logic                     := 'X';             -- reset_n
			avs_s1_write           : in  std_logic                     := 'X';             -- write
			avs_s1_read            : in  std_logic                     := 'X';             -- read
			avs_s1_chipselect      : in  std_logic                     := 'X';             -- chipselect
			avs_s1_byteenable      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			avs_s1_address         : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- address
			avs_s1_writedata       : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			avs_s1_readdata        : out std_logic_vector(15 downto 0)                     -- readdata
		);
	end component mm_bus_counter;

	component CPU_System_cpu_0 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(26 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(26 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component CPU_System_cpu_0;

	component CPU_System_fpga_sdram is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(24 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(12 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component CPU_System_fpga_sdram;

	component CPU_System_jtag_uart_0 is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component CPU_System_jtag_uart_0;

	component CPU_System_onchip_memory2_1 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(12 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component CPU_System_onchip_memory2_1;

	component CPU_System_pio_input_0 is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(7 downto 0)  := (others => 'X')  -- export
		);
	end component CPU_System_pio_input_0;

	component CPU_System_pio_output_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component CPU_System_pio_output_0;

	component CPU_System_pll is
		port (
			refclk   : in  std_logic := 'X'; -- clk
			rst      : in  std_logic := 'X'; -- reset
			outclk_0 : out std_logic;        -- clk
			outclk_1 : out std_logic;        -- clk
			locked   : out std_logic         -- export
		);
	end component CPU_System_pll;

	component CPU_System_sysid is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component CPU_System_sysid;

	component CPU_System_timer_system is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component CPU_System_timer_system;

	component CPU_System_mm_interconnect_0 is
		port (
			pll_outclk0_clk                            : in  std_logic                     := 'X';             -- clk
			cpu_0_reset_reset_bridge_in_reset_reset    : in  std_logic                     := 'X';             -- reset
			cpu_0_data_master_address                  : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			cpu_0_data_master_waitrequest              : out std_logic;                                        -- waitrequest
			cpu_0_data_master_byteenable               : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			cpu_0_data_master_read                     : in  std_logic                     := 'X';             -- read
			cpu_0_data_master_readdata                 : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_0_data_master_write                    : in  std_logic                     := 'X';             -- write
			cpu_0_data_master_writedata                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			cpu_0_data_master_debugaccess              : in  std_logic                     := 'X';             -- debugaccess
			cpu_0_instruction_master_address           : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			cpu_0_instruction_master_waitrequest       : out std_logic;                                        -- waitrequest
			cpu_0_instruction_master_read              : in  std_logic                     := 'X';             -- read
			cpu_0_instruction_master_readdata          : out std_logic_vector(31 downto 0);                    -- readdata
			bridge_component_0_avalon_slave_address    : out std_logic_vector(7 downto 0);                     -- address
			bridge_component_0_avalon_slave_write      : out std_logic;                                        -- write
			bridge_component_0_avalon_slave_read       : out std_logic;                                        -- read
			bridge_component_0_avalon_slave_readdata   : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			bridge_component_0_avalon_slave_writedata  : out std_logic_vector(15 downto 0);                    -- writedata
			bridge_component_0_avalon_slave_byteenable : out std_logic_vector(1 downto 0);                     -- byteenable
			bridge_component_0_avalon_slave_chipselect : out std_logic;                                        -- chipselect
			cpu_0_debug_mem_slave_address              : out std_logic_vector(8 downto 0);                     -- address
			cpu_0_debug_mem_slave_write                : out std_logic;                                        -- write
			cpu_0_debug_mem_slave_read                 : out std_logic;                                        -- read
			cpu_0_debug_mem_slave_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			cpu_0_debug_mem_slave_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			cpu_0_debug_mem_slave_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			cpu_0_debug_mem_slave_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			cpu_0_debug_mem_slave_debugaccess          : out std_logic;                                        -- debugaccess
			fpga_sdram_s1_address                      : out std_logic_vector(24 downto 0);                    -- address
			fpga_sdram_s1_write                        : out std_logic;                                        -- write
			fpga_sdram_s1_read                         : out std_logic;                                        -- read
			fpga_sdram_s1_readdata                     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			fpga_sdram_s1_writedata                    : out std_logic_vector(15 downto 0);                    -- writedata
			fpga_sdram_s1_byteenable                   : out std_logic_vector(1 downto 0);                     -- byteenable
			fpga_sdram_s1_readdatavalid                : in  std_logic                     := 'X';             -- readdatavalid
			fpga_sdram_s1_waitrequest                  : in  std_logic                     := 'X';             -- waitrequest
			fpga_sdram_s1_chipselect                   : out std_logic;                                        -- chipselect
			onchip_memory2_1_s1_address                : out std_logic_vector(12 downto 0);                    -- address
			onchip_memory2_1_s1_write                  : out std_logic;                                        -- write
			onchip_memory2_1_s1_readdata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_memory2_1_s1_writedata              : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_memory2_1_s1_byteenable             : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_memory2_1_s1_chipselect             : out std_logic;                                        -- chipselect
			onchip_memory2_1_s1_clken                  : out std_logic;                                        -- clken
			pio_input_0_s1_address                     : out std_logic_vector(1 downto 0);                     -- address
			pio_input_0_s1_readdata                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_output_0_s1_address                    : out std_logic_vector(1 downto 0);                     -- address
			pio_output_0_s1_write                      : out std_logic;                                        -- write
			pio_output_0_s1_readdata                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_output_0_s1_writedata                  : out std_logic_vector(31 downto 0);                    -- writedata
			pio_output_0_s1_chipselect                 : out std_logic;                                        -- chipselect
			sysid_control_slave_address                : out std_logic_vector(0 downto 0);                     -- address
			sysid_control_slave_readdata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			timer_system_s1_address                    : out std_logic_vector(2 downto 0);                     -- address
			timer_system_s1_write                      : out std_logic;                                        -- write
			timer_system_s1_readdata                   : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			timer_system_s1_writedata                  : out std_logic_vector(15 downto 0);                    -- writedata
			timer_system_s1_chipselect                 : out std_logic;                                        -- chipselect
			timer_timestamp_s1_address                 : out std_logic_vector(2 downto 0);                     -- address
			timer_timestamp_s1_write                   : out std_logic;                                        -- write
			timer_timestamp_s1_readdata                : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			timer_timestamp_s1_writedata               : out std_logic_vector(15 downto 0);                    -- writedata
			timer_timestamp_s1_chipselect              : out std_logic                                         -- chipselect
		);
	end component CPU_System_mm_interconnect_0;

	component CPU_System_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component CPU_System_irq_mapper;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			reset_in1      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal pll_outclk0_clk                                              : std_logic;                     -- pll:outclk_0 -> [bridge_component_0:csi_clockreset_clk, cpu_0:clk, fpga_sdram:clk, irq_mapper:clk, jtag_uart_0:clk, mm_interconnect_0:pll_outclk0_clk, onchip_memory2_1:clk, pio_input_0:clk, pio_output_0:clk, rst_controller:clk, sysid:clock, timer_system:clk, timer_timestamp:clk]
	signal cpu_0_data_master_readdata                                   : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_0_data_master_readdata -> cpu_0:d_readdata
	signal cpu_0_data_master_waitrequest                                : std_logic;                     -- mm_interconnect_0:cpu_0_data_master_waitrequest -> cpu_0:d_waitrequest
	signal cpu_0_data_master_debugaccess                                : std_logic;                     -- cpu_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_0_data_master_debugaccess
	signal cpu_0_data_master_address                                    : std_logic_vector(26 downto 0); -- cpu_0:d_address -> mm_interconnect_0:cpu_0_data_master_address
	signal cpu_0_data_master_byteenable                                 : std_logic_vector(3 downto 0);  -- cpu_0:d_byteenable -> mm_interconnect_0:cpu_0_data_master_byteenable
	signal cpu_0_data_master_read                                       : std_logic;                     -- cpu_0:d_read -> mm_interconnect_0:cpu_0_data_master_read
	signal cpu_0_data_master_write                                      : std_logic;                     -- cpu_0:d_write -> mm_interconnect_0:cpu_0_data_master_write
	signal cpu_0_data_master_writedata                                  : std_logic_vector(31 downto 0); -- cpu_0:d_writedata -> mm_interconnect_0:cpu_0_data_master_writedata
	signal cpu_0_instruction_master_readdata                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_0_instruction_master_readdata -> cpu_0:i_readdata
	signal cpu_0_instruction_master_waitrequest                         : std_logic;                     -- mm_interconnect_0:cpu_0_instruction_master_waitrequest -> cpu_0:i_waitrequest
	signal cpu_0_instruction_master_address                             : std_logic_vector(26 downto 0); -- cpu_0:i_address -> mm_interconnect_0:cpu_0_instruction_master_address
	signal cpu_0_instruction_master_read                                : std_logic;                     -- cpu_0:i_read -> mm_interconnect_0:cpu_0_instruction_master_read
	signal mm_interconnect_0_bridge_component_0_avalon_slave_chipselect : std_logic;                     -- mm_interconnect_0:bridge_component_0_avalon_slave_chipselect -> bridge_component_0:avs_s1_chipselect
	signal mm_interconnect_0_bridge_component_0_avalon_slave_readdata   : std_logic_vector(15 downto 0); -- bridge_component_0:avs_s1_readdata -> mm_interconnect_0:bridge_component_0_avalon_slave_readdata
	signal mm_interconnect_0_bridge_component_0_avalon_slave_address    : std_logic_vector(7 downto 0);  -- mm_interconnect_0:bridge_component_0_avalon_slave_address -> bridge_component_0:avs_s1_address
	signal mm_interconnect_0_bridge_component_0_avalon_slave_read       : std_logic;                     -- mm_interconnect_0:bridge_component_0_avalon_slave_read -> bridge_component_0:avs_s1_read
	signal mm_interconnect_0_bridge_component_0_avalon_slave_byteenable : std_logic_vector(1 downto 0);  -- mm_interconnect_0:bridge_component_0_avalon_slave_byteenable -> bridge_component_0:avs_s1_byteenable
	signal mm_interconnect_0_bridge_component_0_avalon_slave_write      : std_logic;                     -- mm_interconnect_0:bridge_component_0_avalon_slave_write -> bridge_component_0:avs_s1_write
	signal mm_interconnect_0_bridge_component_0_avalon_slave_writedata  : std_logic_vector(15 downto 0); -- mm_interconnect_0:bridge_component_0_avalon_slave_writedata -> bridge_component_0:avs_s1_writedata
	signal mm_interconnect_0_sysid_control_slave_readdata               : std_logic_vector(31 downto 0); -- sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	signal mm_interconnect_0_sysid_control_slave_address                : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sysid_control_slave_address -> sysid:address
	signal mm_interconnect_0_cpu_0_debug_mem_slave_readdata             : std_logic_vector(31 downto 0); -- cpu_0:debug_mem_slave_readdata -> mm_interconnect_0:cpu_0_debug_mem_slave_readdata
	signal mm_interconnect_0_cpu_0_debug_mem_slave_waitrequest          : std_logic;                     -- cpu_0:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_0_debug_mem_slave_waitrequest
	signal mm_interconnect_0_cpu_0_debug_mem_slave_debugaccess          : std_logic;                     -- mm_interconnect_0:cpu_0_debug_mem_slave_debugaccess -> cpu_0:debug_mem_slave_debugaccess
	signal mm_interconnect_0_cpu_0_debug_mem_slave_address              : std_logic_vector(8 downto 0);  -- mm_interconnect_0:cpu_0_debug_mem_slave_address -> cpu_0:debug_mem_slave_address
	signal mm_interconnect_0_cpu_0_debug_mem_slave_read                 : std_logic;                     -- mm_interconnect_0:cpu_0_debug_mem_slave_read -> cpu_0:debug_mem_slave_read
	signal mm_interconnect_0_cpu_0_debug_mem_slave_byteenable           : std_logic_vector(3 downto 0);  -- mm_interconnect_0:cpu_0_debug_mem_slave_byteenable -> cpu_0:debug_mem_slave_byteenable
	signal mm_interconnect_0_cpu_0_debug_mem_slave_write                : std_logic;                     -- mm_interconnect_0:cpu_0_debug_mem_slave_write -> cpu_0:debug_mem_slave_write
	signal mm_interconnect_0_cpu_0_debug_mem_slave_writedata            : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_0_debug_mem_slave_writedata -> cpu_0:debug_mem_slave_writedata
	signal mm_interconnect_0_timer_system_s1_chipselect                 : std_logic;                     -- mm_interconnect_0:timer_system_s1_chipselect -> timer_system:chipselect
	signal mm_interconnect_0_timer_system_s1_readdata                   : std_logic_vector(15 downto 0); -- timer_system:readdata -> mm_interconnect_0:timer_system_s1_readdata
	signal mm_interconnect_0_timer_system_s1_address                    : std_logic_vector(2 downto 0);  -- mm_interconnect_0:timer_system_s1_address -> timer_system:address
	signal mm_interconnect_0_timer_system_s1_write                      : std_logic;                     -- mm_interconnect_0:timer_system_s1_write -> mm_interconnect_0_timer_system_s1_write:in
	signal mm_interconnect_0_timer_system_s1_writedata                  : std_logic_vector(15 downto 0); -- mm_interconnect_0:timer_system_s1_writedata -> timer_system:writedata
	signal mm_interconnect_0_pio_output_0_s1_chipselect                 : std_logic;                     -- mm_interconnect_0:pio_output_0_s1_chipselect -> pio_output_0:chipselect
	signal mm_interconnect_0_pio_output_0_s1_readdata                   : std_logic_vector(31 downto 0); -- pio_output_0:readdata -> mm_interconnect_0:pio_output_0_s1_readdata
	signal mm_interconnect_0_pio_output_0_s1_address                    : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pio_output_0_s1_address -> pio_output_0:address
	signal mm_interconnect_0_pio_output_0_s1_write                      : std_logic;                     -- mm_interconnect_0:pio_output_0_s1_write -> mm_interconnect_0_pio_output_0_s1_write:in
	signal mm_interconnect_0_pio_output_0_s1_writedata                  : std_logic_vector(31 downto 0); -- mm_interconnect_0:pio_output_0_s1_writedata -> pio_output_0:writedata
	signal mm_interconnect_0_pio_input_0_s1_readdata                    : std_logic_vector(31 downto 0); -- pio_input_0:readdata -> mm_interconnect_0:pio_input_0_s1_readdata
	signal mm_interconnect_0_pio_input_0_s1_address                     : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pio_input_0_s1_address -> pio_input_0:address
	signal mm_interconnect_0_timer_timestamp_s1_chipselect              : std_logic;                     -- mm_interconnect_0:timer_timestamp_s1_chipselect -> timer_timestamp:chipselect
	signal mm_interconnect_0_timer_timestamp_s1_readdata                : std_logic_vector(15 downto 0); -- timer_timestamp:readdata -> mm_interconnect_0:timer_timestamp_s1_readdata
	signal mm_interconnect_0_timer_timestamp_s1_address                 : std_logic_vector(2 downto 0);  -- mm_interconnect_0:timer_timestamp_s1_address -> timer_timestamp:address
	signal mm_interconnect_0_timer_timestamp_s1_write                   : std_logic;                     -- mm_interconnect_0:timer_timestamp_s1_write -> mm_interconnect_0_timer_timestamp_s1_write:in
	signal mm_interconnect_0_timer_timestamp_s1_writedata               : std_logic_vector(15 downto 0); -- mm_interconnect_0:timer_timestamp_s1_writedata -> timer_timestamp:writedata
	signal mm_interconnect_0_fpga_sdram_s1_chipselect                   : std_logic;                     -- mm_interconnect_0:fpga_sdram_s1_chipselect -> fpga_sdram:az_cs
	signal mm_interconnect_0_fpga_sdram_s1_readdata                     : std_logic_vector(15 downto 0); -- fpga_sdram:za_data -> mm_interconnect_0:fpga_sdram_s1_readdata
	signal mm_interconnect_0_fpga_sdram_s1_waitrequest                  : std_logic;                     -- fpga_sdram:za_waitrequest -> mm_interconnect_0:fpga_sdram_s1_waitrequest
	signal mm_interconnect_0_fpga_sdram_s1_address                      : std_logic_vector(24 downto 0); -- mm_interconnect_0:fpga_sdram_s1_address -> fpga_sdram:az_addr
	signal mm_interconnect_0_fpga_sdram_s1_read                         : std_logic;                     -- mm_interconnect_0:fpga_sdram_s1_read -> mm_interconnect_0_fpga_sdram_s1_read:in
	signal mm_interconnect_0_fpga_sdram_s1_byteenable                   : std_logic_vector(1 downto 0);  -- mm_interconnect_0:fpga_sdram_s1_byteenable -> mm_interconnect_0_fpga_sdram_s1_byteenable:in
	signal mm_interconnect_0_fpga_sdram_s1_readdatavalid                : std_logic;                     -- fpga_sdram:za_valid -> mm_interconnect_0:fpga_sdram_s1_readdatavalid
	signal mm_interconnect_0_fpga_sdram_s1_write                        : std_logic;                     -- mm_interconnect_0:fpga_sdram_s1_write -> mm_interconnect_0_fpga_sdram_s1_write:in
	signal mm_interconnect_0_fpga_sdram_s1_writedata                    : std_logic_vector(15 downto 0); -- mm_interconnect_0:fpga_sdram_s1_writedata -> fpga_sdram:az_data
	signal mm_interconnect_0_onchip_memory2_1_s1_chipselect             : std_logic;                     -- mm_interconnect_0:onchip_memory2_1_s1_chipselect -> onchip_memory2_1:chipselect
	signal mm_interconnect_0_onchip_memory2_1_s1_readdata               : std_logic_vector(31 downto 0); -- onchip_memory2_1:readdata -> mm_interconnect_0:onchip_memory2_1_s1_readdata
	signal mm_interconnect_0_onchip_memory2_1_s1_address                : std_logic_vector(12 downto 0); -- mm_interconnect_0:onchip_memory2_1_s1_address -> onchip_memory2_1:address
	signal mm_interconnect_0_onchip_memory2_1_s1_byteenable             : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_memory2_1_s1_byteenable -> onchip_memory2_1:byteenable
	signal mm_interconnect_0_onchip_memory2_1_s1_write                  : std_logic;                     -- mm_interconnect_0:onchip_memory2_1_s1_write -> onchip_memory2_1:write
	signal mm_interconnect_0_onchip_memory2_1_s1_writedata              : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_memory2_1_s1_writedata -> onchip_memory2_1:writedata
	signal mm_interconnect_0_onchip_memory2_1_s1_clken                  : std_logic;                     -- mm_interconnect_0:onchip_memory2_1_s1_clken -> onchip_memory2_1:clken
	signal irq_mapper_receiver0_irq                                     : std_logic;                     -- jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                     : std_logic;                     -- timer_system:irq -> irq_mapper:receiver1_irq
	signal irq_mapper_receiver2_irq                                     : std_logic;                     -- timer_timestamp:irq -> irq_mapper:receiver2_irq
	signal cpu_0_irq_irq                                                : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> cpu_0:irq
	signal rst_controller_reset_out_reset                               : std_logic;                     -- rst_controller:reset_out -> [irq_mapper:reset, mm_interconnect_0:cpu_0_reset_reset_bridge_in_reset_reset, onchip_memory2_1:reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                           : std_logic;                     -- rst_controller:reset_req -> [cpu_0:reset_req, onchip_memory2_1:reset_req, rst_translator:reset_req_in]
	signal cpu_0_debug_reset_request_reset                              : std_logic;                     -- cpu_0:debug_reset_request -> rst_controller:reset_in1
	signal reset_reset_n_ports_inv                                      : std_logic;                     -- reset_reset_n:inv -> [pll:rst, rst_controller:reset_in0]
	signal mm_interconnect_0_timer_system_s1_write_ports_inv            : std_logic;                     -- mm_interconnect_0_timer_system_s1_write:inv -> timer_system:write_n
	signal mm_interconnect_0_pio_output_0_s1_write_ports_inv            : std_logic;                     -- mm_interconnect_0_pio_output_0_s1_write:inv -> pio_output_0:write_n
	signal mm_interconnect_0_timer_timestamp_s1_write_ports_inv         : std_logic;                     -- mm_interconnect_0_timer_timestamp_s1_write:inv -> timer_timestamp:write_n
	signal mm_interconnect_0_fpga_sdram_s1_read_ports_inv               : std_logic;                     -- mm_interconnect_0_fpga_sdram_s1_read:inv -> fpga_sdram:az_rd_n
	signal mm_interconnect_0_fpga_sdram_s1_byteenable_ports_inv         : std_logic_vector(1 downto 0);  -- mm_interconnect_0_fpga_sdram_s1_byteenable:inv -> fpga_sdram:az_be_n
	signal mm_interconnect_0_fpga_sdram_s1_write_ports_inv              : std_logic;                     -- mm_interconnect_0_fpga_sdram_s1_write:inv -> fpga_sdram:az_wr_n
	signal rst_controller_reset_out_reset_ports_inv                     : std_logic;                     -- rst_controller_reset_out_reset:inv -> [bridge_component_0:csi_clockreset_reset_n, cpu_0:reset_n, fpga_sdram:reset_n, jtag_uart_0:rst_n, pio_input_0:reset_n, pio_output_0:reset_n, sysid:reset_n, timer_system:reset_n, timer_timestamp:reset_n]

begin

	bridge_component_0 : component mm_bus_counter
		port map (
			csi_clockreset_clk     => pll_outclk0_clk,                                              --       clockreset.clk
			csi_clockreset_reset_n => rst_controller_reset_out_reset_ports_inv,                     -- clockreset_reset.reset_n
			avs_s1_write           => mm_interconnect_0_bridge_component_0_avalon_slave_write,      --     avalon_slave.write
			avs_s1_read            => mm_interconnect_0_bridge_component_0_avalon_slave_read,       --                 .read
			avs_s1_chipselect      => mm_interconnect_0_bridge_component_0_avalon_slave_chipselect, --                 .chipselect
			avs_s1_byteenable      => mm_interconnect_0_bridge_component_0_avalon_slave_byteenable, --                 .byteenable
			avs_s1_address         => mm_interconnect_0_bridge_component_0_avalon_slave_address,    --                 .address
			avs_s1_writedata       => mm_interconnect_0_bridge_component_0_avalon_slave_writedata,  --                 .writedata
			avs_s1_readdata        => mm_interconnect_0_bridge_component_0_avalon_slave_readdata    --                 .readdata
		);

	cpu_0 : component CPU_System_cpu_0
		port map (
			clk                                 => pll_outclk0_clk,                                     --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,            --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                  --                          .reset_req
			d_address                           => cpu_0_data_master_address,                           --               data_master.address
			d_byteenable                        => cpu_0_data_master_byteenable,                        --                          .byteenable
			d_read                              => cpu_0_data_master_read,                              --                          .read
			d_readdata                          => cpu_0_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => cpu_0_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => cpu_0_data_master_write,                             --                          .write
			d_writedata                         => cpu_0_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => cpu_0_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => cpu_0_instruction_master_address,                    --        instruction_master.address
			i_read                              => cpu_0_instruction_master_read,                       --                          .read
			i_readdata                          => cpu_0_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => cpu_0_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => cpu_0_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => cpu_0_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_cpu_0_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_cpu_0_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_cpu_0_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_cpu_0_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_cpu_0_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_cpu_0_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_cpu_0_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_cpu_0_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                 -- custom_instruction_master.readra
		);

	fpga_sdram : component CPU_System_fpga_sdram
		port map (
			clk            => pll_outclk0_clk,                                      --   clk.clk
			reset_n        => rst_controller_reset_out_reset_ports_inv,             -- reset.reset_n
			az_addr        => mm_interconnect_0_fpga_sdram_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_0_fpga_sdram_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_0_fpga_sdram_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_0_fpga_sdram_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_0_fpga_sdram_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_0_fpga_sdram_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_0_fpga_sdram_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_0_fpga_sdram_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_0_fpga_sdram_s1_waitrequest,          --      .waitrequest
			zs_addr        => dram_addr,                                            --  wire.export
			zs_ba          => dram_ba,                                              --      .export
			zs_cas_n       => dram_cas_n,                                           --      .export
			zs_cke         => dram_cke,                                             --      .export
			zs_cs_n        => dram_cs_n,                                            --      .export
			zs_dq          => dram_dq,                                              --      .export
			zs_dqm         => dram_dqm,                                             --      .export
			zs_ras_n       => dram_ras_n,                                           --      .export
			zs_we_n        => dram_we_n                                             --      .export
		);

	jtag_uart_0 : component CPU_System_jtag_uart_0
		port map (
			clk            => pll_outclk0_clk,                           --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,  --             reset.reset_n
			av_chipselect  => jtag_uart_0_avalon_jtag_slave_chipselect,  -- avalon_jtag_slave.chipselect
			av_address     => jtag_uart_0_avalon_jtag_slave_address,     --                  .address
			av_read_n      => jtag_uart_0_avalon_jtag_slave_read_n,      --                  .read_n
			av_readdata    => jtag_uart_0_avalon_jtag_slave_readdata,    --                  .readdata
			av_write_n     => jtag_uart_0_avalon_jtag_slave_write_n,     --                  .write_n
			av_writedata   => jtag_uart_0_avalon_jtag_slave_writedata,   --                  .writedata
			av_waitrequest => jtag_uart_0_avalon_jtag_slave_waitrequest, --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                   --               irq.irq
		);

	onchip_memory2_1 : component CPU_System_onchip_memory2_1
		port map (
			clk        => pll_outclk0_clk,                                  --   clk1.clk
			address    => mm_interconnect_0_onchip_memory2_1_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchip_memory2_1_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchip_memory2_1_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchip_memory2_1_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchip_memory2_1_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchip_memory2_1_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_onchip_memory2_1_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,                   -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,               --       .reset_req
			freeze     => '0'                                               -- (terminated)
		);

	pio_input_0 : component CPU_System_pio_input_0
		port map (
			clk      => pll_outclk0_clk,                           --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,  --               reset.reset_n
			address  => mm_interconnect_0_pio_input_0_s1_address,  --                  s1.address
			readdata => mm_interconnect_0_pio_input_0_s1_readdata, --                    .readdata
			in_port  => in_port_to_the_pio_input_0                 -- external_connection.export
		);

	pio_output_0 : component CPU_System_pio_output_0
		port map (
			clk        => pll_outclk0_clk,                                   --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,          --               reset.reset_n
			address    => mm_interconnect_0_pio_output_0_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pio_output_0_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pio_output_0_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pio_output_0_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pio_output_0_s1_readdata,        --                    .readdata
			out_port   => out_port_from_the_pio_output_0                     -- external_connection.export
		);

	pll : component CPU_System_pll
		port map (
			refclk   => clk_50,                  --  refclk.clk
			rst      => reset_reset_n_ports_inv, --   reset.reset
			outclk_0 => pll_outclk0_clk,         -- outclk0.clk
			outclk_1 => dram_clk_clk,            -- outclk1.clk
			locked   => open                     -- (terminated)
		);

	sysid : component CPU_System_sysid
		port map (
			clock    => pll_outclk0_clk,                                  --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,         --         reset.reset_n
			readdata => mm_interconnect_0_sysid_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_control_slave_address(0)  --              .address
		);

	timer_system : component CPU_System_timer_system
		port map (
			clk        => pll_outclk0_clk,                                   --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,          -- reset.reset_n
			address    => mm_interconnect_0_timer_system_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_timer_system_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_timer_system_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_timer_system_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_timer_system_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver1_irq                           --   irq.irq
		);

	timer_timestamp : component CPU_System_timer_system
		port map (
			clk        => pll_outclk0_clk,                                      --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,             -- reset.reset_n
			address    => mm_interconnect_0_timer_timestamp_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_timer_timestamp_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_timer_timestamp_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_timer_timestamp_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_timer_timestamp_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver2_irq                              --   irq.irq
		);

	mm_interconnect_0 : component CPU_System_mm_interconnect_0
		port map (
			pll_outclk0_clk                            => pll_outclk0_clk,                                              --                       pll_outclk0.clk
			cpu_0_reset_reset_bridge_in_reset_reset    => rst_controller_reset_out_reset,                               -- cpu_0_reset_reset_bridge_in_reset.reset
			cpu_0_data_master_address                  => cpu_0_data_master_address,                                    --                 cpu_0_data_master.address
			cpu_0_data_master_waitrequest              => cpu_0_data_master_waitrequest,                                --                                  .waitrequest
			cpu_0_data_master_byteenable               => cpu_0_data_master_byteenable,                                 --                                  .byteenable
			cpu_0_data_master_read                     => cpu_0_data_master_read,                                       --                                  .read
			cpu_0_data_master_readdata                 => cpu_0_data_master_readdata,                                   --                                  .readdata
			cpu_0_data_master_write                    => cpu_0_data_master_write,                                      --                                  .write
			cpu_0_data_master_writedata                => cpu_0_data_master_writedata,                                  --                                  .writedata
			cpu_0_data_master_debugaccess              => cpu_0_data_master_debugaccess,                                --                                  .debugaccess
			cpu_0_instruction_master_address           => cpu_0_instruction_master_address,                             --          cpu_0_instruction_master.address
			cpu_0_instruction_master_waitrequest       => cpu_0_instruction_master_waitrequest,                         --                                  .waitrequest
			cpu_0_instruction_master_read              => cpu_0_instruction_master_read,                                --                                  .read
			cpu_0_instruction_master_readdata          => cpu_0_instruction_master_readdata,                            --                                  .readdata
			bridge_component_0_avalon_slave_address    => mm_interconnect_0_bridge_component_0_avalon_slave_address,    --   bridge_component_0_avalon_slave.address
			bridge_component_0_avalon_slave_write      => mm_interconnect_0_bridge_component_0_avalon_slave_write,      --                                  .write
			bridge_component_0_avalon_slave_read       => mm_interconnect_0_bridge_component_0_avalon_slave_read,       --                                  .read
			bridge_component_0_avalon_slave_readdata   => mm_interconnect_0_bridge_component_0_avalon_slave_readdata,   --                                  .readdata
			bridge_component_0_avalon_slave_writedata  => mm_interconnect_0_bridge_component_0_avalon_slave_writedata,  --                                  .writedata
			bridge_component_0_avalon_slave_byteenable => mm_interconnect_0_bridge_component_0_avalon_slave_byteenable, --                                  .byteenable
			bridge_component_0_avalon_slave_chipselect => mm_interconnect_0_bridge_component_0_avalon_slave_chipselect, --                                  .chipselect
			cpu_0_debug_mem_slave_address              => mm_interconnect_0_cpu_0_debug_mem_slave_address,              --             cpu_0_debug_mem_slave.address
			cpu_0_debug_mem_slave_write                => mm_interconnect_0_cpu_0_debug_mem_slave_write,                --                                  .write
			cpu_0_debug_mem_slave_read                 => mm_interconnect_0_cpu_0_debug_mem_slave_read,                 --                                  .read
			cpu_0_debug_mem_slave_readdata             => mm_interconnect_0_cpu_0_debug_mem_slave_readdata,             --                                  .readdata
			cpu_0_debug_mem_slave_writedata            => mm_interconnect_0_cpu_0_debug_mem_slave_writedata,            --                                  .writedata
			cpu_0_debug_mem_slave_byteenable           => mm_interconnect_0_cpu_0_debug_mem_slave_byteenable,           --                                  .byteenable
			cpu_0_debug_mem_slave_waitrequest          => mm_interconnect_0_cpu_0_debug_mem_slave_waitrequest,          --                                  .waitrequest
			cpu_0_debug_mem_slave_debugaccess          => mm_interconnect_0_cpu_0_debug_mem_slave_debugaccess,          --                                  .debugaccess
			fpga_sdram_s1_address                      => mm_interconnect_0_fpga_sdram_s1_address,                      --                     fpga_sdram_s1.address
			fpga_sdram_s1_write                        => mm_interconnect_0_fpga_sdram_s1_write,                        --                                  .write
			fpga_sdram_s1_read                         => mm_interconnect_0_fpga_sdram_s1_read,                         --                                  .read
			fpga_sdram_s1_readdata                     => mm_interconnect_0_fpga_sdram_s1_readdata,                     --                                  .readdata
			fpga_sdram_s1_writedata                    => mm_interconnect_0_fpga_sdram_s1_writedata,                    --                                  .writedata
			fpga_sdram_s1_byteenable                   => mm_interconnect_0_fpga_sdram_s1_byteenable,                   --                                  .byteenable
			fpga_sdram_s1_readdatavalid                => mm_interconnect_0_fpga_sdram_s1_readdatavalid,                --                                  .readdatavalid
			fpga_sdram_s1_waitrequest                  => mm_interconnect_0_fpga_sdram_s1_waitrequest,                  --                                  .waitrequest
			fpga_sdram_s1_chipselect                   => mm_interconnect_0_fpga_sdram_s1_chipselect,                   --                                  .chipselect
			onchip_memory2_1_s1_address                => mm_interconnect_0_onchip_memory2_1_s1_address,                --               onchip_memory2_1_s1.address
			onchip_memory2_1_s1_write                  => mm_interconnect_0_onchip_memory2_1_s1_write,                  --                                  .write
			onchip_memory2_1_s1_readdata               => mm_interconnect_0_onchip_memory2_1_s1_readdata,               --                                  .readdata
			onchip_memory2_1_s1_writedata              => mm_interconnect_0_onchip_memory2_1_s1_writedata,              --                                  .writedata
			onchip_memory2_1_s1_byteenable             => mm_interconnect_0_onchip_memory2_1_s1_byteenable,             --                                  .byteenable
			onchip_memory2_1_s1_chipselect             => mm_interconnect_0_onchip_memory2_1_s1_chipselect,             --                                  .chipselect
			onchip_memory2_1_s1_clken                  => mm_interconnect_0_onchip_memory2_1_s1_clken,                  --                                  .clken
			pio_input_0_s1_address                     => mm_interconnect_0_pio_input_0_s1_address,                     --                    pio_input_0_s1.address
			pio_input_0_s1_readdata                    => mm_interconnect_0_pio_input_0_s1_readdata,                    --                                  .readdata
			pio_output_0_s1_address                    => mm_interconnect_0_pio_output_0_s1_address,                    --                   pio_output_0_s1.address
			pio_output_0_s1_write                      => mm_interconnect_0_pio_output_0_s1_write,                      --                                  .write
			pio_output_0_s1_readdata                   => mm_interconnect_0_pio_output_0_s1_readdata,                   --                                  .readdata
			pio_output_0_s1_writedata                  => mm_interconnect_0_pio_output_0_s1_writedata,                  --                                  .writedata
			pio_output_0_s1_chipselect                 => mm_interconnect_0_pio_output_0_s1_chipselect,                 --                                  .chipselect
			sysid_control_slave_address                => mm_interconnect_0_sysid_control_slave_address,                --               sysid_control_slave.address
			sysid_control_slave_readdata               => mm_interconnect_0_sysid_control_slave_readdata,               --                                  .readdata
			timer_system_s1_address                    => mm_interconnect_0_timer_system_s1_address,                    --                   timer_system_s1.address
			timer_system_s1_write                      => mm_interconnect_0_timer_system_s1_write,                      --                                  .write
			timer_system_s1_readdata                   => mm_interconnect_0_timer_system_s1_readdata,                   --                                  .readdata
			timer_system_s1_writedata                  => mm_interconnect_0_timer_system_s1_writedata,                  --                                  .writedata
			timer_system_s1_chipselect                 => mm_interconnect_0_timer_system_s1_chipselect,                 --                                  .chipselect
			timer_timestamp_s1_address                 => mm_interconnect_0_timer_timestamp_s1_address,                 --                timer_timestamp_s1.address
			timer_timestamp_s1_write                   => mm_interconnect_0_timer_timestamp_s1_write,                   --                                  .write
			timer_timestamp_s1_readdata                => mm_interconnect_0_timer_timestamp_s1_readdata,                --                                  .readdata
			timer_timestamp_s1_writedata               => mm_interconnect_0_timer_timestamp_s1_writedata,               --                                  .writedata
			timer_timestamp_s1_chipselect              => mm_interconnect_0_timer_timestamp_s1_chipselect               --                                  .chipselect
		);

	irq_mapper : component CPU_System_irq_mapper
		port map (
			clk           => pll_outclk0_clk,                --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,       -- receiver2.irq
			sender_irq    => cpu_0_irq_irq                   --    sender.irq
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1      => cpu_0_debug_reset_request_reset,    -- reset_in1.reset
			clk            => pll_outclk0_clk,                    --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_timer_system_s1_write_ports_inv <= not mm_interconnect_0_timer_system_s1_write;

	mm_interconnect_0_pio_output_0_s1_write_ports_inv <= not mm_interconnect_0_pio_output_0_s1_write;

	mm_interconnect_0_timer_timestamp_s1_write_ports_inv <= not mm_interconnect_0_timer_timestamp_s1_write;

	mm_interconnect_0_fpga_sdram_s1_read_ports_inv <= not mm_interconnect_0_fpga_sdram_s1_read;

	mm_interconnect_0_fpga_sdram_s1_byteenable_ports_inv <= not mm_interconnect_0_fpga_sdram_s1_byteenable;

	mm_interconnect_0_fpga_sdram_s1_write_ports_inv <= not mm_interconnect_0_fpga_sdram_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of CPU_System
