// CPU_System.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module CPU_System (
		input  wire        clk_50,                         //                    clk_50_clk_in.clk
		output wire [12:0] dram_addr,                      //                             dram.addr
		output wire [1:0]  dram_ba,                        //                                 .ba
		output wire        dram_cas_n,                     //                                 .cas_n
		output wire        dram_cke,                       //                                 .cke
		output wire        dram_cs_n,                      //                                 .cs_n
		inout  wire [15:0] dram_dq,                        //                                 .dq
		output wire [1:0]  dram_dqm,                       //                                 .dqm
		output wire        dram_ras_n,                     //                                 .ras_n
		output wire        dram_we_n,                      //                                 .we_n
		output wire        dram_clk_clk,                   //                         dram_clk.clk
		input  wire [7:0]  in_port_to_the_pio_input_0,     //  pio_input_0_external_connection.export
		output wire [7:0]  out_port_from_the_pio_output_0, // pio_output_0_external_connection.export
		input  wire        reset_reset_n                   //                            reset.reset_n
	);

	wire         pll_outclk0_clk;                                             // pll:outclk_0 -> [cpu_0:clk, fpga_sdram:clk, irq_mapper:clk, jtag_uart_0:clk, mm_interconnect_0:pll_outclk0_clk, onchip_memory2_1:clk, pio_input_0:clk, pio_output_0:clk, rst_controller:clk, sysid:clock, timer_system:clk, timer_timestamp:clk]
	wire  [31:0] cpu_0_data_master_readdata;                                  // mm_interconnect_0:cpu_0_data_master_readdata -> cpu_0:d_readdata
	wire         cpu_0_data_master_waitrequest;                               // mm_interconnect_0:cpu_0_data_master_waitrequest -> cpu_0:d_waitrequest
	wire         cpu_0_data_master_debugaccess;                               // cpu_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_0_data_master_debugaccess
	wire  [26:0] cpu_0_data_master_address;                                   // cpu_0:d_address -> mm_interconnect_0:cpu_0_data_master_address
	wire   [3:0] cpu_0_data_master_byteenable;                                // cpu_0:d_byteenable -> mm_interconnect_0:cpu_0_data_master_byteenable
	wire         cpu_0_data_master_read;                                      // cpu_0:d_read -> mm_interconnect_0:cpu_0_data_master_read
	wire         cpu_0_data_master_write;                                     // cpu_0:d_write -> mm_interconnect_0:cpu_0_data_master_write
	wire  [31:0] cpu_0_data_master_writedata;                                 // cpu_0:d_writedata -> mm_interconnect_0:cpu_0_data_master_writedata
	wire  [31:0] cpu_0_instruction_master_readdata;                           // mm_interconnect_0:cpu_0_instruction_master_readdata -> cpu_0:i_readdata
	wire         cpu_0_instruction_master_waitrequest;                        // mm_interconnect_0:cpu_0_instruction_master_waitrequest -> cpu_0:i_waitrequest
	wire  [26:0] cpu_0_instruction_master_address;                            // cpu_0:i_address -> mm_interconnect_0:cpu_0_instruction_master_address
	wire         cpu_0_instruction_master_read;                               // cpu_0:i_read -> mm_interconnect_0:cpu_0_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_control_slave_readdata;              // sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_control_slave_address;               // mm_interconnect_0:sysid_control_slave_address -> sysid:address
	wire  [31:0] mm_interconnect_0_cpu_0_debug_mem_slave_readdata;            // cpu_0:debug_mem_slave_readdata -> mm_interconnect_0:cpu_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_0_debug_mem_slave_waitrequest;         // cpu_0:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_0_debug_mem_slave_debugaccess;         // mm_interconnect_0:cpu_0_debug_mem_slave_debugaccess -> cpu_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_0_debug_mem_slave_address;             // mm_interconnect_0:cpu_0_debug_mem_slave_address -> cpu_0:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_0_debug_mem_slave_read;                // mm_interconnect_0:cpu_0_debug_mem_slave_read -> cpu_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_0_debug_mem_slave_byteenable;          // mm_interconnect_0:cpu_0_debug_mem_slave_byteenable -> cpu_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_0_debug_mem_slave_write;               // mm_interconnect_0:cpu_0_debug_mem_slave_write -> cpu_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_0_debug_mem_slave_writedata;           // mm_interconnect_0:cpu_0_debug_mem_slave_writedata -> cpu_0:debug_mem_slave_writedata
	wire         mm_interconnect_0_timer_system_s1_chipselect;                // mm_interconnect_0:timer_system_s1_chipselect -> timer_system:chipselect
	wire  [15:0] mm_interconnect_0_timer_system_s1_readdata;                  // timer_system:readdata -> mm_interconnect_0:timer_system_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_system_s1_address;                   // mm_interconnect_0:timer_system_s1_address -> timer_system:address
	wire         mm_interconnect_0_timer_system_s1_write;                     // mm_interconnect_0:timer_system_s1_write -> timer_system:write_n
	wire  [15:0] mm_interconnect_0_timer_system_s1_writedata;                 // mm_interconnect_0:timer_system_s1_writedata -> timer_system:writedata
	wire         mm_interconnect_0_pio_output_0_s1_chipselect;                // mm_interconnect_0:pio_output_0_s1_chipselect -> pio_output_0:chipselect
	wire  [31:0] mm_interconnect_0_pio_output_0_s1_readdata;                  // pio_output_0:readdata -> mm_interconnect_0:pio_output_0_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_output_0_s1_address;                   // mm_interconnect_0:pio_output_0_s1_address -> pio_output_0:address
	wire         mm_interconnect_0_pio_output_0_s1_write;                     // mm_interconnect_0:pio_output_0_s1_write -> pio_output_0:write_n
	wire  [31:0] mm_interconnect_0_pio_output_0_s1_writedata;                 // mm_interconnect_0:pio_output_0_s1_writedata -> pio_output_0:writedata
	wire  [31:0] mm_interconnect_0_pio_input_0_s1_readdata;                   // pio_input_0:readdata -> mm_interconnect_0:pio_input_0_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_input_0_s1_address;                    // mm_interconnect_0:pio_input_0_s1_address -> pio_input_0:address
	wire         mm_interconnect_0_timer_timestamp_s1_chipselect;             // mm_interconnect_0:timer_timestamp_s1_chipselect -> timer_timestamp:chipselect
	wire  [15:0] mm_interconnect_0_timer_timestamp_s1_readdata;               // timer_timestamp:readdata -> mm_interconnect_0:timer_timestamp_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_timestamp_s1_address;                // mm_interconnect_0:timer_timestamp_s1_address -> timer_timestamp:address
	wire         mm_interconnect_0_timer_timestamp_s1_write;                  // mm_interconnect_0:timer_timestamp_s1_write -> timer_timestamp:write_n
	wire  [15:0] mm_interconnect_0_timer_timestamp_s1_writedata;              // mm_interconnect_0:timer_timestamp_s1_writedata -> timer_timestamp:writedata
	wire         mm_interconnect_0_fpga_sdram_s1_chipselect;                  // mm_interconnect_0:fpga_sdram_s1_chipselect -> fpga_sdram:az_cs
	wire  [15:0] mm_interconnect_0_fpga_sdram_s1_readdata;                    // fpga_sdram:za_data -> mm_interconnect_0:fpga_sdram_s1_readdata
	wire         mm_interconnect_0_fpga_sdram_s1_waitrequest;                 // fpga_sdram:za_waitrequest -> mm_interconnect_0:fpga_sdram_s1_waitrequest
	wire  [24:0] mm_interconnect_0_fpga_sdram_s1_address;                     // mm_interconnect_0:fpga_sdram_s1_address -> fpga_sdram:az_addr
	wire         mm_interconnect_0_fpga_sdram_s1_read;                        // mm_interconnect_0:fpga_sdram_s1_read -> fpga_sdram:az_rd_n
	wire   [1:0] mm_interconnect_0_fpga_sdram_s1_byteenable;                  // mm_interconnect_0:fpga_sdram_s1_byteenable -> fpga_sdram:az_be_n
	wire         mm_interconnect_0_fpga_sdram_s1_readdatavalid;               // fpga_sdram:za_valid -> mm_interconnect_0:fpga_sdram_s1_readdatavalid
	wire         mm_interconnect_0_fpga_sdram_s1_write;                       // mm_interconnect_0:fpga_sdram_s1_write -> fpga_sdram:az_wr_n
	wire  [15:0] mm_interconnect_0_fpga_sdram_s1_writedata;                   // mm_interconnect_0:fpga_sdram_s1_writedata -> fpga_sdram:az_data
	wire         mm_interconnect_0_onchip_memory2_1_s1_chipselect;            // mm_interconnect_0:onchip_memory2_1_s1_chipselect -> onchip_memory2_1:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_1_s1_readdata;              // onchip_memory2_1:readdata -> mm_interconnect_0:onchip_memory2_1_s1_readdata
	wire  [12:0] mm_interconnect_0_onchip_memory2_1_s1_address;               // mm_interconnect_0:onchip_memory2_1_s1_address -> onchip_memory2_1:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_1_s1_byteenable;            // mm_interconnect_0:onchip_memory2_1_s1_byteenable -> onchip_memory2_1:byteenable
	wire         mm_interconnect_0_onchip_memory2_1_s1_write;                 // mm_interconnect_0:onchip_memory2_1_s1_write -> onchip_memory2_1:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_1_s1_writedata;             // mm_interconnect_0:onchip_memory2_1_s1_writedata -> onchip_memory2_1:writedata
	wire         mm_interconnect_0_onchip_memory2_1_s1_clken;                 // mm_interconnect_0:onchip_memory2_1_s1_clken -> onchip_memory2_1:clken
	wire         irq_mapper_receiver0_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                    // timer_system:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                    // timer_timestamp:irq -> irq_mapper:receiver2_irq
	wire  [31:0] cpu_0_irq_irq;                                               // irq_mapper:sender_irq -> cpu_0:irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [cpu_0:reset_n, fpga_sdram:reset_n, irq_mapper:reset, jtag_uart_0:rst_n, mm_interconnect_0:cpu_0_reset_reset_bridge_in_reset_reset, onchip_memory2_1:reset, pio_input_0:reset_n, pio_output_0:reset_n, rst_translator:in_reset, sysid:reset_n, timer_system:reset_n, timer_timestamp:reset_n]
	wire         rst_controller_reset_out_reset_req;                          // rst_controller:reset_req -> [cpu_0:reset_req, onchip_memory2_1:reset_req, rst_translator:reset_req_in]
	wire         cpu_0_debug_reset_request_reset;                             // cpu_0:debug_reset_request -> rst_controller:reset_in1

	CPU_System_cpu_0 cpu_0 (
		.clk                                 (pll_outclk0_clk),                                     //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                     //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                  //                          .reset_req
		.d_address                           (cpu_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_0_data_master_read),                              //                          .read
		.d_readdata                          (cpu_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_0_data_master_write),                             //                          .write
		.d_writedata                         (cpu_0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (cpu_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_0_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_0_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (cpu_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (cpu_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                     // custom_instruction_master.readra
	);

	CPU_System_fpga_sdram fpga_sdram (
		.clk            (pll_outclk0_clk),                               //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),               // reset.reset_n
		.az_addr        (mm_interconnect_0_fpga_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_fpga_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_fpga_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_fpga_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_fpga_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_fpga_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_fpga_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_fpga_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_fpga_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (dram_addr),                                     //  wire.export
		.zs_ba          (dram_ba),                                       //      .export
		.zs_cas_n       (dram_cas_n),                                    //      .export
		.zs_cke         (dram_cke),                                      //      .export
		.zs_cs_n        (dram_cs_n),                                     //      .export
		.zs_dq          (dram_dq),                                       //      .export
		.zs_dqm         (dram_dqm),                                      //      .export
		.zs_ras_n       (dram_ras_n),                                    //      .export
		.zs_we_n        (dram_we_n)                                      //      .export
	);

	CPU_System_jtag_uart_0 jtag_uart_0 (
		.clk            (pll_outclk0_clk),                                             //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	CPU_System_onchip_memory2_1 onchip_memory2_1 (
		.clk        (pll_outclk0_clk),                                  //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_1_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_1_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_1_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_1_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_1_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_1_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_1_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),               //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	CPU_System_pio_input_0 pio_input_0 (
		.clk      (pll_outclk0_clk),                           //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_0_pio_input_0_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pio_input_0_s1_readdata), //                    .readdata
		.in_port  (in_port_to_the_pio_input_0)                 // external_connection.export
	);

	CPU_System_pio_output_0 pio_output_0 (
		.clk        (pll_outclk0_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_pio_output_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_output_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_output_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_output_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_output_0_s1_readdata),   //                    .readdata
		.out_port   (out_port_from_the_pio_output_0)                // external_connection.export
	);

	CPU_System_pll pll (
		.refclk   (clk_50),          //  refclk.clk
		.rst      (~reset_reset_n),  //   reset.reset
		.outclk_0 (pll_outclk0_clk), // outclk0.clk
		.outclk_1 (dram_clk_clk),    // outclk1.clk
		.locked   ()                 // (terminated)
	);

	CPU_System_sysid sysid (
		.clock    (pll_outclk0_clk),                                //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_control_slave_address)   //              .address
	);

	CPU_System_timer_system timer_system (
		.clk        (pll_outclk0_clk),                              //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              // reset.reset_n
		.address    (mm_interconnect_0_timer_system_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_system_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_system_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_system_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_system_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                      //   irq.irq
	);

	CPU_System_timer_system timer_timestamp (
		.clk        (pll_outclk0_clk),                                 //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                 // reset.reset_n
		.address    (mm_interconnect_0_timer_timestamp_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_timestamp_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_timestamp_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_timestamp_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_timestamp_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver2_irq)                         //   irq.irq
	);

	CPU_System_mm_interconnect_0 mm_interconnect_0 (
		.pll_outclk0_clk                           (pll_outclk0_clk),                                             //                       pll_outclk0.clk
		.cpu_0_reset_reset_bridge_in_reset_reset   (rst_controller_reset_out_reset),                              // cpu_0_reset_reset_bridge_in_reset.reset
		.cpu_0_data_master_address                 (cpu_0_data_master_address),                                   //                 cpu_0_data_master.address
		.cpu_0_data_master_waitrequest             (cpu_0_data_master_waitrequest),                               //                                  .waitrequest
		.cpu_0_data_master_byteenable              (cpu_0_data_master_byteenable),                                //                                  .byteenable
		.cpu_0_data_master_read                    (cpu_0_data_master_read),                                      //                                  .read
		.cpu_0_data_master_readdata                (cpu_0_data_master_readdata),                                  //                                  .readdata
		.cpu_0_data_master_write                   (cpu_0_data_master_write),                                     //                                  .write
		.cpu_0_data_master_writedata               (cpu_0_data_master_writedata),                                 //                                  .writedata
		.cpu_0_data_master_debugaccess             (cpu_0_data_master_debugaccess),                               //                                  .debugaccess
		.cpu_0_instruction_master_address          (cpu_0_instruction_master_address),                            //          cpu_0_instruction_master.address
		.cpu_0_instruction_master_waitrequest      (cpu_0_instruction_master_waitrequest),                        //                                  .waitrequest
		.cpu_0_instruction_master_read             (cpu_0_instruction_master_read),                               //                                  .read
		.cpu_0_instruction_master_readdata         (cpu_0_instruction_master_readdata),                           //                                  .readdata
		.cpu_0_debug_mem_slave_address             (mm_interconnect_0_cpu_0_debug_mem_slave_address),             //             cpu_0_debug_mem_slave.address
		.cpu_0_debug_mem_slave_write               (mm_interconnect_0_cpu_0_debug_mem_slave_write),               //                                  .write
		.cpu_0_debug_mem_slave_read                (mm_interconnect_0_cpu_0_debug_mem_slave_read),                //                                  .read
		.cpu_0_debug_mem_slave_readdata            (mm_interconnect_0_cpu_0_debug_mem_slave_readdata),            //                                  .readdata
		.cpu_0_debug_mem_slave_writedata           (mm_interconnect_0_cpu_0_debug_mem_slave_writedata),           //                                  .writedata
		.cpu_0_debug_mem_slave_byteenable          (mm_interconnect_0_cpu_0_debug_mem_slave_byteenable),          //                                  .byteenable
		.cpu_0_debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_0_debug_mem_slave_waitrequest),         //                                  .waitrequest
		.cpu_0_debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_0_debug_mem_slave_debugaccess),         //                                  .debugaccess
		.fpga_sdram_s1_address                     (mm_interconnect_0_fpga_sdram_s1_address),                     //                     fpga_sdram_s1.address
		.fpga_sdram_s1_write                       (mm_interconnect_0_fpga_sdram_s1_write),                       //                                  .write
		.fpga_sdram_s1_read                        (mm_interconnect_0_fpga_sdram_s1_read),                        //                                  .read
		.fpga_sdram_s1_readdata                    (mm_interconnect_0_fpga_sdram_s1_readdata),                    //                                  .readdata
		.fpga_sdram_s1_writedata                   (mm_interconnect_0_fpga_sdram_s1_writedata),                   //                                  .writedata
		.fpga_sdram_s1_byteenable                  (mm_interconnect_0_fpga_sdram_s1_byteenable),                  //                                  .byteenable
		.fpga_sdram_s1_readdatavalid               (mm_interconnect_0_fpga_sdram_s1_readdatavalid),               //                                  .readdatavalid
		.fpga_sdram_s1_waitrequest                 (mm_interconnect_0_fpga_sdram_s1_waitrequest),                 //                                  .waitrequest
		.fpga_sdram_s1_chipselect                  (mm_interconnect_0_fpga_sdram_s1_chipselect),                  //                                  .chipselect
		.jtag_uart_0_avalon_jtag_slave_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //     jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                  .write
		.jtag_uart_0_avalon_jtag_slave_read        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                  .read
		.jtag_uart_0_avalon_jtag_slave_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                  .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                  .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                  .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                  .chipselect
		.onchip_memory2_1_s1_address               (mm_interconnect_0_onchip_memory2_1_s1_address),               //               onchip_memory2_1_s1.address
		.onchip_memory2_1_s1_write                 (mm_interconnect_0_onchip_memory2_1_s1_write),                 //                                  .write
		.onchip_memory2_1_s1_readdata              (mm_interconnect_0_onchip_memory2_1_s1_readdata),              //                                  .readdata
		.onchip_memory2_1_s1_writedata             (mm_interconnect_0_onchip_memory2_1_s1_writedata),             //                                  .writedata
		.onchip_memory2_1_s1_byteenable            (mm_interconnect_0_onchip_memory2_1_s1_byteenable),            //                                  .byteenable
		.onchip_memory2_1_s1_chipselect            (mm_interconnect_0_onchip_memory2_1_s1_chipselect),            //                                  .chipselect
		.onchip_memory2_1_s1_clken                 (mm_interconnect_0_onchip_memory2_1_s1_clken),                 //                                  .clken
		.pio_input_0_s1_address                    (mm_interconnect_0_pio_input_0_s1_address),                    //                    pio_input_0_s1.address
		.pio_input_0_s1_readdata                   (mm_interconnect_0_pio_input_0_s1_readdata),                   //                                  .readdata
		.pio_output_0_s1_address                   (mm_interconnect_0_pio_output_0_s1_address),                   //                   pio_output_0_s1.address
		.pio_output_0_s1_write                     (mm_interconnect_0_pio_output_0_s1_write),                     //                                  .write
		.pio_output_0_s1_readdata                  (mm_interconnect_0_pio_output_0_s1_readdata),                  //                                  .readdata
		.pio_output_0_s1_writedata                 (mm_interconnect_0_pio_output_0_s1_writedata),                 //                                  .writedata
		.pio_output_0_s1_chipselect                (mm_interconnect_0_pio_output_0_s1_chipselect),                //                                  .chipselect
		.sysid_control_slave_address               (mm_interconnect_0_sysid_control_slave_address),               //               sysid_control_slave.address
		.sysid_control_slave_readdata              (mm_interconnect_0_sysid_control_slave_readdata),              //                                  .readdata
		.timer_system_s1_address                   (mm_interconnect_0_timer_system_s1_address),                   //                   timer_system_s1.address
		.timer_system_s1_write                     (mm_interconnect_0_timer_system_s1_write),                     //                                  .write
		.timer_system_s1_readdata                  (mm_interconnect_0_timer_system_s1_readdata),                  //                                  .readdata
		.timer_system_s1_writedata                 (mm_interconnect_0_timer_system_s1_writedata),                 //                                  .writedata
		.timer_system_s1_chipselect                (mm_interconnect_0_timer_system_s1_chipselect),                //                                  .chipselect
		.timer_timestamp_s1_address                (mm_interconnect_0_timer_timestamp_s1_address),                //                timer_timestamp_s1.address
		.timer_timestamp_s1_write                  (mm_interconnect_0_timer_timestamp_s1_write),                  //                                  .write
		.timer_timestamp_s1_readdata               (mm_interconnect_0_timer_timestamp_s1_readdata),               //                                  .readdata
		.timer_timestamp_s1_writedata              (mm_interconnect_0_timer_timestamp_s1_writedata),              //                                  .writedata
		.timer_timestamp_s1_chipselect             (mm_interconnect_0_timer_timestamp_s1_chipselect)              //                                  .chipselect
	);

	CPU_System_irq_mapper irq_mapper (
		.clk           (pll_outclk0_clk),                //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.sender_irq    (cpu_0_irq_irq)                   //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_0_debug_reset_request_reset),    // reset_in1.reset
		.clk            (pll_outclk0_clk),                    //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
